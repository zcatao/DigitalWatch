

module watch(
	input clk_1Khz,
	input rst,
	input start,
	input stop,
	input time_out,
	output[23:0] dispbuf
	);
	

endmodule 