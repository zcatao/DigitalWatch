

module disp(
	input[23:0] dispbuf,
	output[23:0] dispout
	);
	
	assign dispout = dispbuf;

endmodule 